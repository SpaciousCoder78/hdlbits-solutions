module top_module( 
    input a, 
    input b, 
    output out );
    xnor xn1(out,a,b);
endmodule
